** Profile: "INA848_Test_Circuit-ina848_transient"  [ H:\OneDrive\Project\Amplifier\simulation\ina848\ina848 test circuit-pspicefiles\ina848_test_circuit\ina848_transient.sim ] 

** Creating circuit file "ina848_transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ina848.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 
.OPTIONS EXPAND
.OPTIONS LIBRARY
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\INA848_Test_Circuit.net" 


.END
